s(R1,p(C1,s(R1,p(C1,R1))))
[100, 1E-6, 100, 1E-6, 100]
[0, 0, 0, 0, 0]
[inf, inf, inf, inf, inf]
