s(R1,p(C1,s(R1,E2)))
[100, 1E-6, 100, 1.5E-6, 0.5]
[0, 0, 0, 0, 0.5]
[inf, inf, inf, inf, 0.5]
