s(C1,p(R1,s(R1,C1)))
[1E-6, 100, 100, 1E-6]
[0, 0, 0, 0]
[inf, inf, inf, inf]
