s(R1,p(C1,s(R1,E2)))
[100, 1E-6, 100, 1.5E-6, 0.85]
[0, 0, 0, 0, 0]
[inf, inf, inf, inf. inf]
