s(p(s(p(s(p(R1,C1),R1),C1),R1),C1),R1)
[100,1e-6,100,1e-6,100,1e-6,100]
[0,0,0,0,0,0,0]
[inf,inf,inf,inf,inf,inf,inf]