s(R1,p(R1,C1),p(R1,C1),p(R1,C1)) % circuit string
[100,100,1e-6,100,1e-6,100,1e-6] % initial parameters
[0,0,0,0,0,0,0] % lower boundary conditions
[inf,inf,inf,inf,inf,inf,inf] % upper boundary conditions
