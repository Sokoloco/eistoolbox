s(R1,p(R1,E2)
[100, 100, 1E-6, 0.85]
[0, 0, 0, 0]
[inf, inf, inf, inf]
