s(R1,p(R1,E2))
[240, 3000, 1.5E-6, 0.85]
[0, 0, 0, 0]
[inf, inf, inf, inf]
