s(R1,p(R1,C1),p(R1,C1),p(R1,C1))
[100,100,1e-6,100,1e-6,100,1e-6]
[0,0,0,0,0,0,0]
[inf,inf,inf,inf,inf,inf,inf]
