s(R1,p(s(R1,E2),C1))
[100, 100, 1E-6, 0.5, 1E-6]
[0, 0, 0, 0.5, 0]
[inf, inf, inf, 0.5, inf]
