s(R1,p(R1,C1))
[240, 3000, 1.5E-6]
[0, 0, 0]
[inf, inf, inf]
% randles cell