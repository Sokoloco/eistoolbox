s(R1,p(R1,C1))
[100, 100, 1E-6]
[0, 0, 0]
[inf, inf, inf]
